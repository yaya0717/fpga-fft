module divider #(
	parameter		A_LEN = 8,
	parameter		B_LEN = 4)(
	input								CLK,						// ʱ���ź�
	input								RSTN,                // ��λ�źţ�����Ч
	input								EN,                  // ����������Ч,ʹ���ź�
	input [A_LEN-1:0]				Dividend,				//������
	input	[B_LEN-1:0]				Divisor,					//����
	
	output [A_LEN-1:0]			Quotient,				//��
	output [B_LEN-1:0]			Mod,						//��
	output							RDY);
	
	wire [A_LEN-1:0]				Quotient_reg		[A_LEN-1:0];
	wire [B_LEN-1:0] 				Mod_reg				[A_LEN-1:0];
	wire [A_LEN-1:0]				Dividend_ini_reg	[A_LEN-1:0];
	wire [A_LEN-1:0]				rdy;
	wire [B_LEN-1:0]				Divisor_reg			[A_LEN-1:0];
	
	// ��ʼ����һ��Div_cellģ�飬��������ı������ͳ���
	Div_cell	#(.A_LEN(A_LEN),.B_LEN(B_LEN))	Divider(
		.CLK(CLK),
		.RSTN(RSTN),
		.EN(EN),
		.Dividend({{(B_LEN){1'b0}}, Dividend[A_LEN-1]}),		// �������������λ��0ƴ��
		.Divisor(Divisor),	
		.Dividend_i(Dividend),
		.Quotient_i('b0),
 
		.Quotient(Quotient_reg[A_LEN-1]),
		.Mod(Mod_reg[A_LEN-1]),		
		.Dividend_o(Dividend_ini_reg[A_LEN-1]),
		.Divisor_o(Divisor_reg[A_LEN-1]),
		.RDY(rdy[A_LEN-1])
		);
	
	// ���ɶ��Div_cellģ�飬������ˮ�߼���ṹ
	genvar i;
	
	generate 
		for(i=A_LEN-2;i>=0;i=i-1) begin : Div_flow_loop
			Div_cell	#(.A_LEN(A_LEN),.B_LEN(B_LEN))	Divider(
				.CLK(CLK),
				.RSTN(RSTN),
				.EN(rdy[i+1]),
				.Dividend({Mod_reg[i+1], Dividend_ini_reg[i+1][i]}),	// ��ǰ��������һ��������λƴ��
				.Divisor(Divisor_reg[i+1]),	
				.Dividend_i(Dividend_ini_reg[i+1]),
				.Quotient_i(Quotient_reg[i+1]),
		
				.Quotient(Quotient_reg[i]),
				.Mod(Mod_reg[i]),		
				.Dividend_o(Dividend_ini_reg[i]),
				.Divisor_o(Divisor_reg[i]),
				.RDY(rdy[i])
				);	
		end
	endgenerate
	
	assign RDY=rdy[0];
	assign Quotient = Quotient_reg[0];
	assign Mod = Mod_reg[0]; 
	
endmodule
 
 
module Div_cell#(
	parameter						A_LEN = 8,
	parameter						B_LEN = 4
	)(
	input											CLK,						// ʱ���ź�
	input											RSTN,						// ��λ�źţ�����Ч
	input											EN,						// ����������Ч,ʹ���ź�
	input [B_LEN:0]							Dividend,				//������,����һ�����ݵ����������ⲿģ��ƴ�ӵ�ԭʼ����������һλ
	input	[B_LEN-1:0]							Divisor,					//��һ�����ݵĳ���
	input [A_LEN-1:0]							Dividend_i,				//ԭʼ������
	input [A_LEN-1:0]							Quotient_i,				//��һ�����ݵ���
	
	output reg [A_LEN-1:0]					Quotient,				//��,���ݵ���һ��
	output reg [B_LEN-1:0]					Mod,						//��,Ҳ����һ���ı�����
	output reg [A_LEN-1:0]					Dividend_o,				//ԭʼ������
	output reg [B_LEN-1:0]					Divisor_o,				//ԭʼ����								
	output reg									RDY);
	
	always @(posedge CLK or negedge RSTN) begin
		if(!RSTN) begin													// �첽��λ���������мĴ���
			Quotient <=	'b0;
			Mod <= 'b0;	
			Dividend_o <= 'b0;
			Divisor_o <= 'b0;
			RDY <= 'b0;	
		end else if(EN) begin											// ��ʹ���ź���Чʱ�����г�������
			RDY <= 1'b1;
			Dividend_o <= Dividend_i;
			Divisor_o <= Divisor;
			if(Dividend>={1'b0,Divisor}) begin						// ��ǰ���������ڵ��ڳ���ʱ���̼�1����������
				Quotient <= (Quotient_i<<1)+1'b1;
				Mod <= Dividend-{1'b0,Divisor};
			end else begin																
				Quotient <= (Quotient_i<<1)+1'b0;					// ��ǰ������С�ڳ���ʱ���̲��䣬��������
				Mod <= Dividend;
			end
		end else begin														// ��ʹ���ź���Чʱ���������мĴ���
			Quotient <=	'b0;
			Mod <= 'b0;	
			Dividend_o <= 'b0;
			Divisor_o <= 'b0;
			RDY <= 'b0;
		end
	end
	
endmodule