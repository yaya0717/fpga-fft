module encoder(
                clk, 
                rst_n,
                A, //A��
                B, //B��
                left,
                right
);

input   clk,rst_n;
input   A,B;
output left,right;
reg [3:0] testcnt;

//10ms������������������
reg ok_10ms;
reg [31:0]cnt0;
always@(posedge clk,negedge rst_n)
begin
    if(!rst_n)begin
        cnt0 <= 0;
        ok_10ms <= 1'b0;
    end
    else begin
        if(cnt0 < 32'd5_9999)begin
            cnt0 <= cnt0 + 1'b1;
            ok_10ms <= 1'b0;
        end
        else begin
            cnt0 <= 0;
            ok_10ms <= 1'b1;
        end
    end
end


//ͬ��/���� A��B
reg A_reg,A_reg0;
reg B_reg,B_reg0;
wire A_Debounce;
wire B_Debounce;
always@(posedge clk,negedge rst_n)begin
    if(!rst_n)begin
        A_reg <= 1'b1;
        A_reg0 <= 1'b1;
        B_reg <= 1'b1;
        B_reg0 <= 1'b1;
    end
    else begin
        if(ok_10ms)begin
            A_reg <= A;
            A_reg0 <= A_reg;
            B_reg <= B;
            B_reg0 <= B_reg;
        end
    end
end

assign A_Debounce = A_reg0 && A_reg && A;
assign B_Debounce = B_reg0 && B_reg && B;


//���������A���������أ��½��ؼ�⡣
reg A_Debounce_reg;
wire A_posedge,A_negedge;
always@(posedge clk,negedge rst_n)begin
    if(!rst_n)begin
        A_Debounce_reg <= 1'b1;
    end
    else begin
        A_Debounce_reg <= A_Debounce;
    end
end
assign A_posedge = !A_Debounce_reg && A_Debounce;
assign A_negedge = A_Debounce_reg && !A_Debounce;


//��AB�����������Ϊ��������
reg rotary_right;
reg rotary_left;
always@(posedge clk,negedge rst_n)begin
    if(!rst_n)begin
        rotary_right <= 1'b1;
        rotary_left <= 1'b1;
    end
    else begin
        //A��������ʱ�����BΪ�͵�ƽ������ת����������ת
        if(A_posedge && !B_Debounce)begin
            rotary_right <= 1'b1;
        end
        //A������ʱ�����BΪ�ߵ�ƽ������ת����������ת
        else if(A_posedge && B_Debounce)begin
            rotary_left <= 1'b1;
        end
        //A���½���BΪ�ߵ�ƽ����һ����ת����
        else if(A_negedge && B_Debounce)begin
            rotary_right <= 1'b0;
        end
        //A���½���BΪ�͵�ƽ����һ����ת����
        else if(A_negedge && !B_Debounce)begin
            rotary_left <= 1'b0;
        end
    end
end


//ͨ����������������Է��֣�
//"rotary_right"Ϊ�����ص�ʱ���־��һ����ת
//"rotary_left" Ϊ�����ص�ʱ���־��һ����ת
//���´����Ƕ�����������ؼ��
reg rotary_right_reg,rotary_left_reg;
wire rotary_right_pos,rotary_left_pos;
always@(posedge clk,negedge rst_n)begin
    if(!rst_n)begin
        rotary_right_reg <= 1'b1;
        rotary_left_reg <= 1'b1;
    end
    else begin
        rotary_right_reg <= rotary_right;
        rotary_left_reg <= rotary_left;
    end
end

assign rotary_right_pos = !rotary_right_reg && rotary_right;
assign rotary_left_pos = !rotary_left_reg && rotary_left;

//���ڲ��Եļ����� ��ת+1 ��ת-1
always@(posedge clk,negedge rst_n)begin
    if(!rst_n)
         testcnt <= 4'd0;
    else if(rotary_right_pos)
         testcnt <= testcnt + 4'd1;
    else if(rotary_left_pos)
         testcnt <= testcnt - 4'd1;
end

assign right = rotary_right_pos;
assign left = rotary_left_pos;

endmodule